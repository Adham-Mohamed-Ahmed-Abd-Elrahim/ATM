module rom #(parameter ROM_DATA_WIDTH = 17,
                       ROM_MEM_SIZE   = 64)
(
    // input & output ports
	input  wire                             clk,
	input  wire                             read_enable,
	input  wire  [$clog2(ROM_MEM_SIZE)-1:0] address,
	output wire  [ROM_DATA_WIDTH-1:0]       data_out
);

(*rom_style = "block" *) reg [ROM_DATA_WIDTH-1:0] data; // to infer block ram Resources

//-----------------------------------------------------------
//----------------------- Memory Logic ----------------------
//-----------------------------------------------------------
always  @(posedge clk) begin

    if(read_enable) begin

        case (address)

			'd0:  data <= 'b1000010000100011_1;		'd1:  data <= 'b0001100001000111_1;
			'd2:  data <= 'b0100001001001001_1;		'd3:  data <= 'b0001001100011001_0;
			'd4:  data <= 'b0101100100010111_0;		'd5:  data <= 'b1000000101100101_1;
			'd6:  data <= 'b0001010001100000_1;		'd7:  data <= 'b0010011010011000_1;
			'd8:  data <= 'b0100001010001001_1;		'd9:  data <= 'b0011000110011000_1;
			'd10: data <= 'b1000000101010101_1;		'd11: data <= 'b0100000101101000_1;
			'd12: data <= 'b0110011101001001_1;		'd13: data <= 'b0101010001000000_1;
			'd14: data <= 'b0110001001010001_1;		'd15: data <= 'b1001010001010011_0;
			'd16: data <= 'b1001010010010001_0;		'd17: data <= 'b0010000000000101_1;
			'd18: data <= 'b1000010110010001_1;		'd19: data <= 'b0100000100010100_1;
			'd20: data <= 'b0001100100000111_1;		'd21: data <= 'b0100010001010000_1;
			'd22: data <= 'b0101010110010011_1;		'd23: data <= 'b1001011001001001_0;
			'd24: data <= 'b0100001101000011_1;		'd25: data <= 'b0001000100010001_1;
			'd26: data <= 'b1000011100110111_1;		'd27: data <= 'b0001100110011001_1;
			'd28: data <= 'b0101001100000101_0;		'd29: data <= 'b1000011001001001_1;
			'd30: data <= 'b0101011000110010_1;		'd31: data <= 'b0101000000011001_1;
			'd32: data <= 'b1000001000000100_1;		'd33: data <= 'b0001000110000011_1;
			'd34: data <= 'b0110000101010011_1;		'd35: data <= 'b0100011100000010_1;
			'd36: data <= 'b1001100001100110_1;		'd37: data <= 'b1000001000010010_1;
			'd38: data <= 'b0001010010000101_1;		'd39: data <= 'b0010011100010100_1;
			'd40: data <= 'b0101000001110001_1;		'd41: data <= 'b0111001100100110_1;
			'd42: data <= 'b0011100110001000_1;		'd43: data <= 'b0100001000111001_1;
			'd44: data <= 'b1001001010010011_1;		'd45: data <= 'b1001010110000010_1;
			'd46: data <= 'b0100011001101001_1;		'd47: data <= 'b1001000010000111_1;
			'd48: data <= 'b0011100101110010_1;		'd49: data <= 'b0001011101000100_1;
			'd50: data <= 'b0101011101000000_1;		'd51: data <= 'b0110100101000111_0;
			'd52: data <= 'b1001000000110110_0;		'd53: data <= 'b1001011010000110_1;
			'd54: data <= 'b0111100100101001_1;		'd55: data <= 'b0111100000110001_1;
			'd56: data <= 'b0111001110010000_1;		'd57: data <= 'b0111001100010011_1;
			'd58: data <= 'b0111100100000101_1;		'd59: data <= 'b1001011101101001_1;
			'd60: data <= 'b0100001101100011_1;		'd61: data <= 'b0001011101000111_1;
			'd62: data <= 'b0011000101010110_1;		'd63: data <= 'b0010100110010011_1;

        endcase
    end
end

assign data_out = data;

endmodule