
int i=0;
int k=0;
integer user_count=0;
integer operation_count=0;
int cancel_first = 1;
task maintask;
  $display("============================================================");
  $display("=====================main task=====================",$realtime);
  $display("============================================================");
 fork  
  begin 
    clock_gen();
  end
  begin
    reset_init();

		
      card_rand();
  end
/*begin
  check_idle();
end*/
 join_any 
endtask //automatic

//--------------------------------------------------
task clock_gen;
  $display("============================================================");
  $display("=====================clock_gen =====================",$realtime);
  $display("============================================================");
while(1) begin
clk=0;
#(clk_period/2);
clk=1;
#(clk_period/2);
cover_states.sample();
cover_states_trans.sample();
cg_op_choice_inst.sample();
cg_input_card_pin_inst.sample();

toggle_1.sample();
toggle_2.sample();
toggle_3.sample();
//toggle_4.sample();
toggle_trans_en_int.sample();
toggle_5.sample();
toggle_6.sample();
toggle_7.sample();
//toggle_8.sample();
toggle_valid_inst.sample();
toggle_9.sample();
toggle_10.sample();
toggle_wren_inst.sample();

end
endtask 
//---------------------------------------------------
task reset_init;
  $display("============================================================");
  $display("=====================reset =====================",$realtime);
  $display("============================================================");

rst_n=1;
#12ns;
rst_n=0;
#12ns;
rst_n=1;
atm_init='0;
enter=0;
cancel=0;
//language_choice=0;
endtask 

task static card_rand();
  $display("============================================================");
  $display("===================== card_rand  =====================",$realtime);
  $display("============================================================");
  //initializing atm_capacity
  atm_capacity=$urandom % 10000000  ;
  pulse(atm_init);
  repeat(1000)begin
 // Card Insertion 
    user_count=user_count+1;
  input_card_pin=$urandom % (DEPTH);   //// Randomize 
  pulse(insert);
  check_card(valid_card_out);
   if( cancel_en==1'b1 || card_spell_out ||password_rand || (valid_card_out==1'b0)) continue;
  //if(valid_card_out);
	begin// language choice
  language_choice=$urandom % 2;  //randomized
	pulse(enter);
	// operation_choice
  repeat(5)begin
    operation_count=operation_count+1;
    operation_rand();
    @(posedge clk);
    if(atm_top_inst.atm_inst.current_state==IDLE)break;
  end
  pulse(cancel);
  @(posedge clk);
  operation_count=0;
	/*repeat(10)begin
	if(atm_top_inst.atm_inst.current_state==IDLE)
	begin
	break;
	end
	else
	operation_rand();
	end*/
	/*// operation_choice
	op_choice=op;
	pulse(enter);*/
	end
    end
  
  
  endtask

task static operation_rand();
  $display("============================================================");
  $display("===================== operation_rand  =====================",$realtime);
  $display("============================================================");
  operation_choice_rand=  $urandom % (4);
  op_choice=operation_choice_rand;
  pulse(enter);
  //pulse(enter);  
  case(operation_choice_rand)
    WITHDRAWAL_OP:begin 
     //  cancel_rand(); //cancel_Randomization
       withdrawal_val_set();
       cancel_rand(); //cancel_Randomization
    //   @(posedge clk);
      // $display("cancel=%d , abort=%d , cancel_en=%d ,card_spell_out=%d ",done,abort,cancel_en,card_spell_out);
       if((done==1'b1) || abort==1'b1 || cancel_en==1'b1 || card_spell_out==1'b1);
    end
 TRANSFER_OP:begin
  transfer_val_set();   
  cancel_rand(); //cancel_Randomization

  if((done==1'b1)|| (abort==1'b1) || cancel_en==1'b1);
 end
BALANCE_SERVICE_OP:begin
  $display("============================================================");
  $display("===================== BALANCE_SERVICE_OP  =====================",$realtime);
  $display("============================================================");
  @(posedge(done));
end
DEPOSITE_OP:begin
  $display("============================================================");
  $display("===================== DEPOSITE_OP  =====================",$realtime);
  $display("============================================================"); 
  deposite_val_set();
  cancel_rand(); //cancel_Randomization
@(posedge(done));
  //if(done==1'b1 || (cancel_en && atm_top_inst.atm_inst.timer_en_r==1'b0) ) ;
 end
  endcase 
 
    // To set value to be withdrew

endtask 
//---------------------------------------------------
 task automatic pulse(ref logic  signal);
  @(posedge clk) begin
    signal=1'b1;
  end
  @(posedge clk) begin
    signal=1'b0;
  end
endtask

task check_card( output bit valid_card);
  $display("============================================================");
  $display("===================== check_card  =====================",$realtime);
  $display("============================================================");
  cancel_rand(); //cancel_Randomization
  if(cancel_en!=1'b1)begin
  password_rand=$urandom %2; //password_randomization
  //input_password=rom[pin_card][]+$urand(1);
   input_password=rom[input_card_pin][ROM_DATA_WIDTH-1:1]+password_rand; 
   pulse(enter);
  $display("ref_password=%d",rom[input_card_pin][ROM_DATA_WIDTH-1:1], "input_password=%d",input_password);
  //check_password
if((input_password==rom[input_card_pin][ROM_DATA_WIDTH-1:1])&& rom[input_card_pin][0]==1'b1)begin
valid_card=1'b1;
end
else 
begin 
  valid_card=1'b0;
end
 end
  
endtask 
//--------------------------------------------------
/*
task seq_generator(logic [OP_CHOICE_SIZE-1:0] op);
  $display("============================================================");
  $display("===================== seq_generator  =====================",$realtime);
  $display("============================================================");

  //initializing atm_capacity
  atm_capacity=$urandom % 10000000  ;
  pulse(atm_init);
// Card Insertion 
  input_card_pin=$urandom % (DEPTH);   //// Randomize 
  //$display();
 // input_card_pin=0;
  pulse(insert);
  check_card(valid_card_out);
  if(valid_card_out);
begin// language choice
language_choice=1'b1; //English
pulse(enter);
// operation_choice
op_choice=op;
pulse(enter);
end
//seq_generator(op);
  //check_idle();
//cancel_rand(); //cancel_Randomization
endtask 
*/


task transfer_val_set();
  $display("============================================================");
  $display("===================== transfer_val_set  =====================",$realtime);
  $display("============================================================");
  //initializing withdrawal value
  transfer_value=$urandom %(32767);
  transfer_card_pin=1;
  $display("trnasfer_value=%d",withdrawal_value);
  pulse(enter);
  pulse(enter);
endtask 

task withdrawal_val_set();
  $display("============================================================");
  $display("===================== withdrawal_val_set  =====================",$realtime);
  $display("============================================================");
  //initializing withdrawal value
  if(cancel_first) begin
    pulse(cancel);
    cancel_first = 0;
  end
  withdrawal_value=$urandom %(32767);
  $display("Withdrawal_value=%d",withdrawal_value);
  pulse(enter);
  pulse(enter);
endtask 
task deposite_val_set();
  $display("============================================================");
  $display("===================== deposite_val_set  =====================",$realtime);
  $display("============================================================");
  //initializing withdrawal value
  deposite_value=$urandom %(32767);
  $display("deposite_value_value=%d",withdrawal_value);
  pulse(enter);
 pulse(enter);
endtask 

task cancel_rand();
cancel_en=$urandom % 2;
if(cancel_en)begin
  pulse(cancel);
end
endtask

task cancel_rand_cond();
output logic cancel_en;
cancel_en=$urandom % 2;
if(cancel_en)begin
  pulse(cancel);
end
endtask

task check_idle(logic [OP_CHOICE_SIZE-1:0] op);
//while(1)begin
if(atm_top_inst.atm_inst.current_state==IDLE)begin
 //repeat(5) @(posedge clk);
//seq_generator(op);
end
endtask
//----------------------------------------------
